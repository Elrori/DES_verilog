/**************************************************************************************
*   Name        :des_pc2.v
*   Description :DES subkeys pc2,part of des_top.v 
*                输入最高位编号1，最低为编号64,其他类似
*   Origin      :20181228
*   Author      :helrori2011@gmail.com
**************************************************************************************/
module des_pc2
(
    input   wire [1:28] li_28,
    input   wire [1:28] ri_28,
    output  wire [1:48] kout_48
);
wire [1:56]in_56;
assign in_56 = {li_28,ri_28};
assign kout_48 = {
in_56[14], in_56[17], in_56[11], in_56[24], in_56[1],  in_56[5], 
in_56[3],  in_56[28], in_56[15], in_56[6],  in_56[21], in_56[10],
in_56[23], in_56[19], in_56[12], in_56[4],  in_56[26], in_56[8], 
in_56[16], in_56[7],  in_56[27], in_56[20], in_56[13], in_56[2],

in_56[41], in_56[52], in_56[31], in_56[37], in_56[47], in_56[55], 
in_56[30], in_56[40], in_56[51], in_56[45], in_56[33], in_56[48], 
in_56[44], in_56[49], in_56[39], in_56[56], in_56[34], in_56[53], 
in_56[46], in_56[42], in_56[50], in_56[36], in_56[29], in_56[32]

};
endmodule